module DIO(input clk,rstn,
            input [15:0] d,
            input pre,
            input bs,
            input nxt,
            output [7:0] an,
            output [6:0] seg
);

//对输入去抖动并同步化
wire DS_bs,DS_pre,DS_nxt;
wire [15:0] DS_d;
wire [3:0] En_d;

reg [15:0] DR;
reg [4:0] AR;
reg [15:0] DReg;
reg [15:0] DNxt;

reg [7:0] Count;

reg [4:0] wa;

reg [15:0] wd;

reg we;
wire [15:0] RD;

reg [2:0] CS,NS;

reg [1:0] T;   // {nxt,pre}

parameter s0 = 3'b000,s1 = 3'b001,s2 = 3'b010,s3 = 3'b011,s4 = 3'b100,s5 = 3'b101;


deSyn desyn_bs(clk,rstn,bs,DS_bs);
deSyn desyn_pre(clk,rstn,pre,DS_pre);
deSyn desyn_nxt(clk,rstn,nxt,DS_nxt);

deSyn desyn_d0(clk,rstn,d[0],DS_d[0]);
deSyn desyn_d1(clk,rstn,d[1],DS_d[1]);
deSyn desyn_d2(clk,rstn,d[2],DS_d[2]);
deSyn desyn_d3(clk,rstn,d[3],DS_d[3]);
deSyn desyn_d4(clk,rstn,d[4],DS_d[4]);
deSyn desyn_d5(clk,rstn,d[5],DS_d[5]);
deSyn desyn_d6(clk,rstn,d[6],DS_d[6]);
deSyn desyn_d7(clk,rstn,d[7],DS_d[7]);
deSyn desyn_d8(clk,rstn,d[8],DS_d[8]);
deSyn desyn_d9(clk,rstn,d[9],DS_d[9]);
deSyn desyn_d10(clk,rstn,d[10],DS_d[10]);
deSyn desyn_d11(clk,rstn,d[11],DS_d[11]);
deSyn desyn_d12(clk,rstn,d[12],DS_d[12]);
deSyn desyn_d13(clk,rstn,d[13],DS_d[13]);
deSyn desyn_d14(clk,rstn,d[14],DS_d[14]);
deSyn desyn_d15(clk,rstn,d[15],DS_d[15]);




encode ECD(DNxt,En_d);

register_file RF(.clk(clk),.ra0(AR),.rd0(RD),.wa(AR),.wd(DR),.we(we));

dynimage DIS(clk,rstn,Count,DR,an,seg);

always @(posedge clk,negedge rstn) begin
    if(!rstn) 
        CS <= s0;
    else CS <= NS;
    
end

/*
s0:默认状态
s1:读出数字并显示
s2:输入数字
s3:保存数字
s4:退格
s5:显示上一个数字或下一个数字
*/

always @(*) begin
    case(CS)
    s0: NS = s1;
    s1: NS = s2;
    s2: begin
      if(T[1]||T[0])  NS = s5;
      else if(DS_bs) NS = s4;
      else if(DNxt) NS = s3;
      else NS = s2;
    end
    s3: NS = s2;
    s4: NS = s2;
    s5: NS = s1;  
    endcase      
end


always @(posedge clk,negedge rstn) begin
    if(!rstn) begin
      DNxt <= 0;
      DReg <= 0;
      AR <= 0;
      DR <= 0;
      Count <= 0;
      we <= 0;
    end
    else begin
      DNxt <= DS_d - DReg;
      DReg <= DS_d;
      case(NS)
      s1:begin
          DR <= RD;
          we <= 0;
      end
      s2:begin
         T <= {DS_nxt,DS_pre};
         we <= 0;
      end 
      s3:begin
          DR <= (DR<<4)+En_d;
          we <= 1;
      end 
      s4:begin
         DR <=  DR >> 4;
         we <= 1;
      end 
      s5:begin
         we = 0;
        if(T[1]) begin
          AR <= AR +1;
          Count <= Count +1;
        end 
        if(T[0]) begin
          AR <= AR -1;
          Count <= Count -1;
        end 
      end 
      endcase
    end
end

endmodule










//其他模块

module deSyn(input clk,rstn,input x,output y);
wire de_x;
debounce DB(clk,rstn,x,de_x);
Synchron SYN(de_x,clk,rstn,y);
endmodule

module debounce(input clk,rstn,               
                input x,
                output reg y);
parameter  Cnt0 = 3'b000, Cnt1 = 3'b001,Assign0 = 3'b010,Assign1=3'b011,Default = 3'b111;   //刚开始进入默认状态，两个计数状态，两个赋值状态    
reg [2:0] CS,NS;
reg [19:0] Count;
reg y_reg;
always @(posedge clk,negedge rstn) begin          //异步复位
    if(!rstn)begin
      CS <= Default;
      y_reg <= 0;
    end 
    else begin
      CS <= NS;
    y_reg <= y;
    end 
end

always @(posedge clk,negedge rstn) begin
  if(!rstn) Count <=0;
  else begin
    case(CS)
       Default: Count <= 0;
    Cnt0 :begin
      Count <= Count+1;
    end 
    Cnt1: Count <= Count+1;
    Assign0: Count <= 0;
    Assign1: Count <= 0;

  endcase
  end

  
end

always @(*) begin
    y = y_reg;
    NS = Default;
    case (CS) 
    Default: begin
      y = 0;
      if(x == 1) NS = Cnt1;
      else NS = Cnt0;
    end
    Cnt0:begin
       if(Count == 100000) begin
         NS = Assign0;
       end 
       else if(x == 0)begin
         NS = Cnt0;
       end    
       else begin
         NS = Default;
       end      
    end
    Cnt1:begin
       if(Count == 100000) begin
         NS = Assign1;
       end 
       else if(x == 1)begin
         NS = Cnt1;
       end    
       else begin
         NS = Default;
       end      
    end
    Assign0: begin
           y = 0;
      if(x == 0)
        NS = Assign0;                
      else 
         NS = Default;              //只有极个别才在此刻为1
    end
    Assign1:begin
      y = 1;
      if(x == 1) NS = Assign1;
      else NS = Default;                  //只有极个别才在此刻为1
    end
    endcase
end
endmodule





module Synchron(input x,input clk,rstn,
                output y);
reg s1,s2;
reg s;

always @(posedge clk) begin
    if(~rstn ) begin
      s1 <= 0;
      s2 <= 0;
      s <= 0;
    end
    else begin
      s1 <= x;
      s2 <= s1;
      s <= s2;
    end
end
assign y = (!s)&s2;
endmodule





module  register_file # (
    parameter AW = 5,		//地址宽度
    parameter DW = 16		//数据宽度
)(
    input clk,			//时钟
    input [AW-1:0] ra0, ra1,		//读地址
    output [DW-1:0] rd0, rd1,	//读数据
    input [AW-1:0] wa, 		//写地址
    input [DW-1:0] wd,		//写数据
    input we			//写使能
);
    reg [DW-1:0] rf [0: (1<<AW)-1];		//寄存器堆
    assign rd0 = rf[ra0], rd1 = rf[ra1];	//读操作
    
    always  @ (posedge  clk)
        if (we)  rf[wa]  <=  wd;		//写操作
endmodule

module encode(input [15:0] In,output reg [3:0] Out );
    always @(*) begin
        case(In)
        16'b0000_0000_0000_0001: Out = 4'b0000;
        16'b0000_0000_0000_0010: Out = 4'b0001;
        16'b0000_0000_0000_0100: Out = 4'b0010;
        16'b0000_0000_0000_1000: Out = 4'b0011;
        16'b0000_0000_0001_0000: Out = 4'b0100;
        16'b0000_0000_0010_0000: Out = 4'b0101;
        16'b0000_0000_0100_0000: Out = 4'b0110;
        16'b0000_0000_1000_0000: Out = 4'b0111;
        16'b0000_0001_0000_0000: Out = 4'b1000;
        16'b0000_0010_0000_0000: Out = 4'b1001;
        16'b0000_0100_0000_0000: Out = 4'b1010;
        16'b0000_1000_0000_0000: Out = 4'b1011;
        16'b0001_0000_0000_0000: Out = 4'b1100;
        16'b0010_0000_0000_0000: Out = 4'b1101;
        16'b0100_0000_0000_0000: Out = 4'b1110;
        16'b1000_0000_0000_0000: Out = 4'b1111;
        endcase       
    end

endmodule

module dynimage(
                input clk,rstn,
                input [7:0] Cnt,
                input [15:0] d,
                output reg [7:0] an,
                output reg [6:0] seg);

                wire clkd;        //分频时钟
                reg [3:0] DIn;
                wire [6:0] DOut;
        frequdivision  FreDivClk(clk,~rstn,clkd);
        Decoder7Seg decoder(DIn,DOut);

parameter s0 = 3'b000, s1 = 3'b001,s2 = 3'b010,s3 = 3'b011,s4 = 3'b100,s5 = 3'b101;
reg [2:0] CS,NS;


always @(posedge clkd,negedge rstn) begin  //异步初始化
    if(~rstn) CS <= s0;
    else CS <= NS;
end

always @(*) begin
      case(CS)
      s0 : begin 
          DIn = d[3:0];  
          an = 8'b1111_1110;
          seg = DOut; 
          NS = s1;
      end
      s1 : begin
        DIn = d[7:4];
        seg = DOut;
        NS = s2;
        an = 8'b1111_1101;
      end
      s2 : begin
        DIn = d[11:8];
        seg = DOut;
        NS = s3;
        an = 8'b1111_1011;  
        
      end
      s3 : begin
        DIn = d[15:12];
        seg = DOut;
        NS = s4;
        an = 8'b1111_0111;
      end
      s4 :begin
        DIn = Cnt[3:0];
        seg = DOut;
        NS = s5;
        an = 8'b1011_1111;
      end
      s5 :begin
        DIn = Cnt[7:4];
        seg = DOut;
        NS = s0;
        an = 8'b0111_1111;
      end
      endcase
end
    

endmodule





module frequdivision #(parameter N = 200000,RST_VLU = 0)(input clk,rst, 
output reg out);  //分频器 N = 100000 ~ 2000000
reg [19:0] cnt ;
always @(posedge clk) begin
   if(rst)  cnt <= RST_VLU;
   else if(cnt == (N-1)) cnt <= 0;
   else cnt <= cnt + 1;
end
always @(posedge clk) begin
    if(rst) out <= 0;
    else if(cnt == (N-2)) out <= 1;
    else out <= 0;
end
endmodule

module Decoder7Seg(            //7段译码管
input wire [3:0] In,
output reg [6:0] Out
    );
always @ (*)
    begin
    case(In)
        4'b0000: Out = 7'b000_0001;
        4'b0001: Out = 7'b100_1111;
        4'b0010: Out = 7'b001_0010;
        4'b0011: Out = 7'b000_0110;
        4'b0100: Out = 7'b100_1100;
        4'b0101: Out = 7'b010_0100;
        4'b0110: Out = 7'b010_0000;
        4'b0111: Out = 7'b000_1111;
        4'b1000: Out = 7'b000_0000;
        4'b1001: Out = 7'b000_0100;
        4'b1010: Out = 7'b000_1000;  //A
        4'b1011: Out = 7'b110_0000;  //b
        4'b1100: Out = 7'b011_0001;  //C
        4'b1101: Out = 7'b100_0010;  //d
        4'b1110: Out = 7'b011_0000;  //E
        4'b1111: Out = 7'b011_1000;  //F
    endcase
    end       
endmodule